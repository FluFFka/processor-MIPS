`ifndef __FUNCT_VH
`define __FUNCT_VH

`define FUNCT_ADD   6'b100000
`define FUNCT_ADDU  6'b100001
`define FUNCT_SUB   6'b100010
`define FUNCT_SUBU  6'b100011
`define FUNCT_SLT   6'b101010
`define FUNCT_SLTU  6'b101011

`endif // __FUNCT_VH
